typedef enum bit {WRITE = 1'b0, READ = 1'b1} i2c_op_t;

parameter int I2C_DATA_WIDTH = 8;
parameter int I2C_ADDR_WIDTH = 7;
