class i2cmb_generator_compulsory_test extends ncsu_component;




endclass
