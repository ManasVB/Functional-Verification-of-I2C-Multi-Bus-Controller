    Mac OS X            	   2   �      �                                      ATTR       �   �   <                  �   <  com.apple.quarantine q/0081;5c328d63;Chrome;B223B03D-48DA-4FE1-9C4C-13E4708B682F 