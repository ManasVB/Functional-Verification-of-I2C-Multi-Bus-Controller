parameter int WB_DATA_WIDTH = 8;
parameter int WB_ADDR_WIDTH = 2;
