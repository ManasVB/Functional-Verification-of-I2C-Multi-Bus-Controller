class i2cmb_dut_functionality_test extends ncsu_component;


endclass
