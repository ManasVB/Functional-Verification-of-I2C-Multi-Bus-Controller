parameter int WB_DATA_WIDTH = 8;
parameter int WB_ADDR_WIDTH = 2;

parameter CSR_Reg = 8'h00;
parameter DPR_Reg = 8'h01;
parameter CMDR_Reg = 8'h02;
parameter FSMR_Reg = 8'h03;
