class i2cmb_register_test extends ncsu_component;


endclass
